library verilog;
use verilog.vl_types.all;
entity AdderControl is
    port(
        CLOCK_50        : in     vl_logic
    );
end AdderControl;
